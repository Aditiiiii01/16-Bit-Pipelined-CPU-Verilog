module ex_mem(
    input clk,
    input reset,
    input [15:0] alu_result_in,
    input [15:0] reg_data2_in,   // for store instructions
    input [3:0] rd_in,
    input reg_write_in,
    input mem_read_in,
    input mem_write_in,
    output reg [15:0] alu_result_out,
    output reg [15:0] reg_data2_out,
    output reg [3:0] rd_out,
    output reg reg_write_out,
    output reg mem_read_out,
    output reg mem_write_out
);

always @(posedge clk or posedge reset) begin
    if (reset) begin
        alu_result_out <= 16'b0;
        reg_data2_out <= 16'b0;
        rd_out <= 4'b0;
        reg_write_out <= 0;
        mem_read_out <= 0;
        mem_write_out <= 0;
    end else begin
        alu_result_out <= alu_result_in;
        reg_data2_out <= reg_data2_in;
        rd_out <= rd_in;
        reg_write_out <= reg_write_in;
        mem_read_out <= mem_read_in;
        mem_write_out <= mem_write_in;
    end
end

endmodule
